LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY processor IS
    PORT(
        clk       : IN std_logic;
        reset     : IN std_logic;
        -- I/O Ports
        IN_PORT   : IN std_logic_vector(31 downto 0);
        OUT_PORT  : OUT std_logic_vector(31 downto 0);

        -- Interrupt signals
        INTR_IN   : IN std_logic;

        -- debugging
        PC_debug       : OUT std_logic_vector(31 downto 0);
        instruction_debug : OUT std_logic_vector(31 downto 0);
        ALU_result_debug : OUT std_logic_vector(31 downto 0);
        CCR_debug       : OUT std_logic_vector(2 downto 0)
    );
END processor;

ARCHITECTURE processor_arch OF processor IS

    -- Constants
    constant RESET_VECTOR : std_logic_vector(31 downto 0) := x"00000000";
    constant INTR_VECTOR  : std_logic_vector(31 downto 0) := x"00000004";

    -- IF Stage Signals
    signal PC_value, PC_plus_4, next_PC : std_logic_vector(31 downto 0);
    signal instruction, PC_branch_addr : std_logic_vector(31 downto 0);
    signal PC_stall, PC_write_enable : std_logic;

    -- IF/ID Pipeline Register Signals
    signal IF_ID_Inst, IF_ID_PCPlus4, IF_ID_IN_PORT : std_logic_vector(31 downto 0);
    signal IF_ID_Write, IF_ID_Flush : std_logic;

    -- ID Stage Signals
    signal opcode : std_logic_vector(6 downto 0);
    signal Rsrc1,Rdst,Rsrc2 : std_logic_vector(2 downto 0);
    signal imm_16bit : std_logic_vector(15 downto 0);

    -- Control Unit Signals
    signal Raddr_Sel, RTI_sig, Branch_sig : std_logic;
    signal Int_Jump_Sel, ALU_A, ALU_B, CCR_En : std_logic;
    signal Int_Idx, J_Type : std_logic_vector(1 downto 0);
    signal ALU_Op : std_logic_vector(2 downto 0);
    signal Mem_Write_En, Mem_Read_En, Stack_En, PCsrc : std_logic;
    signal Stack_Inc,Stack_Dec,  Mem_Op : std_logic;
    signal Mem_Addr_Sel, Mem_Write_Sel : std_logic_vector(1 downto 0);
    signal WE1, WE2, OUT_En, HLT_sig : std_logic;
    signal WB_Wadrr_Sel : std_logic_vector(1 downto 0);
    signal WB_Wdata_Sel : std_logic_vector(2 downto 0);

    -- Register File Signals
    signal Reg_Rdata1, Reg_Rdata2 : std_logic_vector(31 downto 0);  -- 32-bit from register file
    signal Rdata1_32bit, Rdata2_32bit : std_logic_vector(31 downto 0);  -- 32-bit converted
    signal Reg_WE1, Reg_WE2 : std_logic;
    signal Reg_Waddr1, Reg_Waddr2 : std_logic_vector(2 downto 0);
    signal Reg_Wdata1, Reg_Wdata2 : std_logic_vector(31 downto 0);

    -- Mux for Raddr1 selection (based on Raddr_Sel)
    signal Raddr1_selected : std_logic_vector(2 downto 0);
    
    signal CCR_in, CCR_out_sig : std_logic_vector(2 downto 0);
    signal PC_we, SP_we, CCR_we : std_logic;
    
    -- Sign Extender Signals
    signal imm_extended, offset_extended : std_logic_vector(31 downto 0);

    -- Hazard Detection Signals
    signal control_mux, insert_nop : std_logic;

    -- ID/EX Pipeline Register Signals
    signal ID_EX_CCR_En, ID_EX_RTI, ID_EX_Int_Jump, ID_EX_Branch : std_logic;
    signal ID_EX_Int_Idx, ID_EX_J_Type : std_logic_vector(1 downto 0);
    signal ID_EX_Mem_Write_En, ID_EX_Mem_Read_En, ID_EX_Stack_En : std_logic;
    signal ID_EX_PCsrc, ID_EX_Stack_Inc,ID_EX_Stack_Dec ,ID_EX_Mem_Op, ID_EX_ALU_A, ID_EX_ALU_B : std_logic;
    signal ID_EX_ALU_Op : std_logic_vector(2 downto 0);
    signal ID_EX_WE1, ID_EX_WE2, ID_EX_OUT_En : std_logic;
    signal ID_EX_WB_Wadrr_Sel : std_logic_vector(1 downto 0);
    signal ID_EX_WB_Wdata_Sel : std_logic_vector(2 downto 0);
    signal ID_EX_PCPlus4, ID_EX_Rdata1, ID_EX_Rdata2 : std_logic_vector(31 downto 0);
    signal ID_EX_Rsrc1, ID_EX_Rsrc2, ID_EX_Rdst : std_logic_vector(2 downto 0);
    signal ID_EX_imm, ID_EX_offset : std_logic_vector(31 downto 0);
    signal ID_EX_IN_PORT : std_logic_vector(31 downto 0);
    signal ID_EX_Wdata_Sel: STD_LOGIC_VECTOR(2 downto 0);
    signal ID_EX_Waddr_Sel: STD_LOGIC_VECTOR(1 downto 0);


    signal ID_EX_Mem_Addr_Sel : STD_LOGIC_VECTOR(1 downto 0);
    signal ID_EX_Mem_Wdata_Sel : STD_LOGIC_VECTOR(1 downto 0);
    -- EX Stage Signals
    signal ALU_op1, ALU_op2, ALU_result : std_logic_vector(31 downto 0);
    signal CCR_updated, CCR_reserved_sig, CCR_OUT : std_logic_vector(2 downto 0);
    signal EX_CCR_En : std_logic;
    signal EX_RTI, Flags_saved: std_logic;
    signal branch_taken, jump_target_sel : std_logic;
    signal jump_target : std_logic_vector(31 downto 0);
    signal Int_Address, Final_Branch_Adrr : std_logic_vector(31 downto 0);

    -- Forwarding Signals
    signal ForwardA, ForwardB : std_logic_vector(1 downto 0);
    signal EX_MEM_RegWrite, MEM_WB_RegWrite : std_logic;

    -- EX/MEM Pipeline Register Signals
    signal EX_MEM_Mem_Write_En, EX_MEM_Mem_Read_En, EX_MEM_Stack_En,EX_MEM_Stack_Dec : std_logic;
    signal EX_MEM_PCsrc, EX_MEM_WE1, EX_MEM_WE2, EX_MEM_OUT_En, EX_MEM_Stack_Inc : std_logic;
    signal EX_MEM_ALU_result, EX_MEM_Rdata1, EX_MEM_Rdata2 : std_logic_vector(31 downto 0);
    signal EX_MEM_Rdst, EX_MEM_Rsrc1, EX_MEM_Rsrc2 : std_logic_vector(2 downto 0);
    signal EX_MEM_imm : std_logic_vector(31 downto 0);
    signal EX_MEM_PCPlus4 : std_logic_vector(31 downto 0);
    signal EX_MEM_BR_ADDR : std_logic_vector(31 downto 0);
    signal EX_MEM_Waddr_Sel: STD_LOGIC_VECTOR(1 downto 0);
    signal EX_MEM_Wdata_Sel: STD_LOGIC_VECTOR(2 downto 0);
    signal EX_MEM_Mem_Op : STD_LOGIC;
    signal EX_MEM_Mem_Addr_Sel : STD_LOGIC_VECTOR(1 downto 0);
    signal EX_MEM_Mem_Wdata_Sel : STD_LOGIC_VECTOR(1 downto 0);

    -- MEM Stage Signals
    signal Mem_Addr, Mem_Write_Data, Mem_Read_Data : std_logic_vector(31 downto 0);
    signal SP_value, SP_next : std_logic_vector(31 downto 0);
    signal SP_enable, SP_load : std_logic;

    -- MEM/WB Pipeline Register Signals
    signal MEM_WB_WE1, MEM_WB_WE2, MEM_WB_OUT_En : std_logic;
    signal MEM_WB_ALU_result, MEM_WB_Mem_Data, MEM_WB_Rdata1 : std_logic_vector(31 downto 0);
    signal MEM_WB_Rdst,MEM_WB_Rsrc1,MEM_WB_Rsrc2 : std_logic_vector(2 downto 0);
    signal MEM_WB_imm : std_logic_vector(31 downto 0);
    signal MEM_WB_IN_PORT : std_logic_vector(31 downto 0);
    signal MEM_WB_Wdata_Sel : std_logic_vector(2 downto 0);
    signal MEM_WB_Waddr_Sel : std_logic_vector(1 downto 0);


    -- WB Stage Signals
    signal WB_Write_Data, WB_Write_Addr : std_logic_vector(31 downto 0);
    signal WB_WE, WB_WE2_sig : std_logic;

BEGIN

    -- ====== INSTRUCTION FETCH ======
    -- PC
    PC_Unit_inst: entity work.PC_Unit
        Port Map(
            clk => clk,
            reset => reset,
            stall => PC_stall,
            PCSrc => PCsrc,
            M0 => RESET_VECTOR,
            PC_out => PC_value,
            PC_branch => EX_MEM_BR_ADDR
        );

    PC_debug <= PC_value;

    -- Memory
    Memory_inst: entity work.Memory
        Port Map(
            clk => clk,
            reset=>  reset,
            Mem_write => EX_MEM_Mem_Write_En,
            Mem_Read => EX_MEM_Mem_Read_En,
            Mem_Addr => Mem_Addr,
            Write_data => Mem_Write_Data,
            Read_data => Mem_Read_Data
        );

    instruction_debug <= IF_ID_Inst;

    -- ====== IF/ID REGISTER ======

    F_D_Register_inst: entity work.F_D_Register
        Port Map(
            CLK => clk,
            RST => reset,
            EN => IF_ID_Write,
            CLR => IF_ID_Flush,
            Inst => Mem_Read_Data,
            PCPlus4 => PC_value,
            IN_Port => IN_PORT,
            Inst_Out => IF_ID_Inst,
            PCPlus4_Out => IF_ID_PCPlus4,
            IN_Out => IF_ID_IN_PORT
        );

    -- ====== STAGE 2: INSTRUCTION DECODE ======

    -- Instruction
    opcode <= IF_ID_Inst(6 downto 0);
    Rsrc1 <= IF_ID_Inst(9 downto 7);
    Rsrc2 <= IF_ID_Inst(12 downto 10);
    Rdst <= IF_ID_Inst(15 downto 13);
    imm_16bit <= IF_ID_Inst(31 downto 16);

    -- Control Unit
    Control_Unit_inst: entity work.Control_Unit
        Port Map(
            opcode => opcode,
            HW_INT => INTR_IN,
            SW_INT => IF_ID_Inst(16),
            Raddr_Sel => Raddr_Sel,
            RTI => RTI_sig,
            Branch => Branch_sig,
            Int_Jump_Sel => Int_Jump_Sel,
            Int_Idx => Int_Idx,
            J_Type => J_Type,
            ALU_A => ALU_A,
            ALU_B => ALU_B,
            ALU_Op => ALU_Op,
            CCR_En => CCR_En,
            Mem_Write_En => Mem_Write_En,
            Mem_Read_En => Mem_Read_En,
            Stack_En => Stack_En,
            PCsrc => PCsrc,
            Stack_Inc => Stack_Inc,
            Mem_Op => Mem_Op,
            Mem_Addr_Sel => Mem_Addr_Sel,
            Mem_Write_Sel => Mem_Write_Sel,
            WE1 => WE1,
            WE2 => WE2,
            WB_Wadrr_Sel => WB_Wadrr_Sel,
            OUT_En => OUT_En,
            WB_Wdata_Sel => WB_Wdata_Sel,
            HLT => HLT_sig
        );

    -- 1. Mux for Raddr1 selection (Raddr_Sel)
    -- 0: Read from Rsrc1, 1: Read from Rdst
    -- not, inc, out, in , push ,pop, ldm
    Raddr1_selected <= Rdst when opcode = "0011100" or opcode = "0011110" or opcode = "0001110" or opcode = "0001010" or  opcode = "0001001" or opcode = "1000101" or opcode = "1001100" else Rsrc1;

    -- 2. Register File with correct connections
    Register_file_inst: entity work.Register_file
        Port Map(
            clk => clk,
            rst => reset,
            WE1 => Reg_WE1,
            WE2 => Reg_WE2,
            Raddr1 => Raddr1_selected,
            Raddr2 => Rsrc2,
            Waddr1 => Reg_Waddr1,
            Waddr2 => Reg_Waddr2,
            Wdata1 => Reg_Wdata1,
            Wdata2 => Reg_Wdata2,
            Rdata1 => Reg_Rdata1,
            Rdata2 => Reg_Rdata2
        );


    CCR_debug <= CCR_in;

    -- Sign Extenders
    Sign_Extender_imm: entity work.Sign_Extender
        Port Map(
            imm_in => imm_16bit,
            imm_out => imm_extended
        );

    --  Hazard Detection Unit
    Hazard_Detection_Unit_inst: entity work.Hazard_Detection_Unit
        Port Map(
            ID_EX_MemRead => ID_EX_Mem_Read_En,
            ID_EX_Rdst => ID_EX_Rdst,
            IF_ID_Rsrc1 => Rsrc1,
            IF_ID_Rsrc2 => Rsrc2,
            Branch => Branch_sig,
            Jump => PCsrc,
            Mem_Op => EX_MEM_Mem_Op,
            PC_Write => PC_write_enable,
            IF_ID_Write => IF_ID_Write,
            Control_Mux => control_mux,
            IF_ID_CLR => IF_ID_Flush
        );

    PC_stall <= not PC_write_enable;
    insert_nop <= control_mux;

    -- ====== ID/EX REGISTER ======

    D_E_Register_inst: entity work.D_E_Register
        Port Map(
            CLK => clk,
            RST => reset,
            EN => '1',
            CLR => insert_nop,
            CCR_EN => CCR_En,
            RTI => RTI_sig,
            INT_Jump => Int_Jump_Sel,
            INT_IDX => Int_Idx,
            MEM_W => Mem_Write_En,
            Branch => Branch_sig,
            Mem_Wdata_Sel => Mem_Write_Sel,
            MemRead => Mem_Read_En,
            J_Type => J_Type,
            MEM_OP => Mem_Op,
            MEM_SEL => Mem_Addr_Sel,
            OUT_EN => OUT_En,
            ALU_A => ALU_A,
            ALUOp => ALU_Op,
            WE1 => WE1,
            WE2 => WE2,
            MEM_R => '0',
            PCSRC => PCsrc,
            PCPlus4 => IF_ID_PCPlus4,
            Rdata1 => Reg_Rdata1,
            Rdata2 => Reg_Rdata2,
            Raddr1 => Raddr1_selected,
            Raddr2 => Rsrc2,
            Rdst => Rdst,
            Imm => imm_extended,
            IN_Port => IF_ID_IN_PORT,
            ALU_B => ALU_B,
            WB_Wdata_Sel => WB_Wdata_Sel,
            WB_Waddr_Sel => WB_Wadrr_Sel,
            Stack_en => Stack_En,
            Stack_inc => Stack_Inc,
            Stack_dec => Stack_Dec,
            CCR_EN_Out => ID_EX_CCR_En,
            RTI_Out => ID_EX_RTI,
            INT_Jump_Out => ID_EX_Int_Jump,
            INT_IDX_Out => ID_EX_Int_Idx,
            MEM_W_Out => ID_EX_Mem_Write_En,
            Branch_Out => ID_EX_Branch,
            Mem_Wdata_Sel_Out => ID_EX_Mem_Wdata_Sel,
            MemRead_Out => ID_EX_Mem_Read_En,
            J_Type_Out => ID_EX_J_Type,
            MEM_OP_Out => ID_EX_Mem_Op,
            MEM_SEL_Out => ID_EX_Mem_Addr_Sel,
            OUT_EN_Out => ID_EX_OUT_En,
            ALU_A_Out => ID_EX_ALU_A,
            ALUOp_Out => ID_EX_ALU_Op,
            WE1_Out => ID_EX_WE1,
            WE2_Out => ID_EX_WE2,
            MEM_R_Out => open,
            PCSRC_Out => ID_EX_PCsrc,
            Stack_en_Out => ID_EX_Stack_En,
            Stack_Inc_Out => ID_EX_Stack_Inc,
            Stack_Dec_Out => ID_EX_Stack_Dec,
            PCPlus4_Out => ID_EX_PCPlus4,
            Rdata1_Out => ID_EX_Rdata1,
            Rdata2_Out => ID_EX_Rdata2,
            Raddr1_Out => ID_EX_Rsrc1,
            Raddr2_Out => ID_EX_Rsrc2,
            Rdst_Out => ID_EX_Rdst,
            Imm_Out => ID_EX_imm,
            IN_Out => ID_EX_IN_PORT,
            ALU_B_Out => ID_EX_ALU_B,
            WB_Waddr_Sel_Out => ID_EX_Waddr_Sel,
            WB_Wdata_Sel_Out => ID_EX_Wdata_Sel
        );

    -- ====== EXECUTE ======

    -- 4. Forwarding Unit with Rsrc1 and Rsrc2
    Forwarding_Unit_inst: entity work.Forward_unit
        Port Map(
            EX_MEM_RegWrite => EX_MEM_WE1,
            MEM_WB_RegWrite => MEM_WB_WE1,
            EX_MEM_Rdst => EX_MEM_Rdst,
            MEM_WB_Rdst => MEM_WB_Rdst,
            ID_EX_Rsrc1 => ID_EX_Rsrc1,
            ID_EX_Rsrc2 => ID_EX_Rsrc2,
            ForwardA => ForwardA,
            ForwardB => ForwardB
        );

    -- ALU  Mux (Forwarding)
    process(ForwardA, ForwardB, ID_EX_Rdata1, ID_EX_Rdata2,
            EX_MEM_ALU_result, MEM_WB_ALU_result, ID_EX_ALU_B, ID_EX_imm)
    begin
        -- ALU Operand A (rsrc1)
        case ForwardA is
            when "00" => ALU_op1 <= ID_EX_Rdata1;
            when "01" => ALU_op1 <= EX_MEM_ALU_result;
            when "10" => ALU_op1 <= MEM_WB_ALU_result;
            when others => ALU_op1 <= ID_EX_Rdata1;
        end case;

        -- ALU Operand B (rsrc2 or immediate)
        if ID_EX_ALU_B = '1' then
            -- Use immediate
            ALU_op2 <= std_logic_vector(resize(signed(ID_EX_imm), 32));
        else
            -- Use Rsrc2
            case ForwardB is
                when "00" => ALU_op2 <= ID_EX_Rdata2;
                when "01" => ALU_op2 <= EX_MEM_ALU_result;
                when "10" => ALU_op2 <= MEM_WB_ALU_result;
                when others => ALU_op2 <= ID_EX_Rdata2;
            end case;
        end if;
    end process;

    -- ALU
    ALU_inst: entity work.ALU
        Port Map
        (
            op1 => ALU_op1,
            op2 => ALU_op2,
            alu_op => ID_EX_ALU_Op, 
           
            alu_out => ALU_result,
            ccr_out =>  CCR_OUT,
            ccr_update => CCR_updated
        );
    
        
    ALU_result_debug <= ALU_result;

    -- CCR update
    --CCR_we <= ID_EX_CCR_En;
    
    CCR_TOP_inst: entity work.CCR_Top
        port map
        (
            clk             => clk,
            reset           => reset,
            ccr_en          => ccr_en,
            int_j           => ID_EX_Int_Jump,
            RTI             => ID_EX_RTI,
            alu_ccr         => CCR_OUT,
            ccr_update      => CCR_updated,
            ccr_out         => CCR_in
        );
    --CCR_in <= "111";
    -- Conditional Branch MUX
    process(ID_EX_J_Type, CCR_in, ID_EX_imm, ID_EX_PCPlus4)
    begin
        branch_taken <= '0';
        jump_target <= (others => '0');

        case ID_EX_J_Type is
            when "00" =>  -- JZ
                branch_taken <= CCR_in(0) and ID_EX_Branch;
            when "01" =>  -- JN
                branch_taken <= CCR_in(1) and ID_EX_Branch;
            when "10" =>  -- JC
                branch_taken <= CCR_in(2) and ID_EX_Branch;
            when "11" =>  -- JMP
                branch_taken <= '1';
            when others =>
                branch_taken <= '0';
        end case;
    end process;

    -- Interrupt address mux
    Int_Address <= x"0000000" & "00" & ID_EX_Int_Idx;

    -- Interrupt/Imm address selection
    jump_target <= ID_EX_imm(31 downto 2) & "00" when ID_EX_Int_Jump = '0' else Int_Address;
    Final_Branch_Adrr <= ID_EX_PCPlus4 when branch_taken = '0' else jump_target;

    -- ====== EX/MEM REGISTER ======

    E_M_Register_inst: entity work.E_M_Register
        Port Map(
            CLK => clk,
            RST => reset,
            EN => '1',
            MemRead => ID_EX_Mem_Read_En,
            MEM_OP => ID_EX_Mem_Op,
            MEM_SEL => ID_EX_Mem_Addr_Sel,
            MEM_R => '0',
            ALURes => ALU_result,
            Raddr1 => ID_EX_Rsrc1,
            Raddr2 => ID_EX_Rsrc2,
            Rdst => ID_EX_Rdst,
            Rdata1 => ALU_op1,
            Rdata2 => ALU_op2,
            Mem_Wdata_Sel => ID_EX_Mem_Wdata_Sel,
            WE1 => ID_EX_WE1,
            WE2 => ID_EX_WE2,
            IN_Port => '0',
            PCSRC => ID_EX_PCsrc,
            Stack_En => ID_EX_Stack_En,
            Stack_Inc => ID_EX_Stack_Inc,
            Stack_Dec => ID_EX_Stack_Dec,
            BR_ADDR => jump_target,
            MEM_W => ID_EX_Mem_Write_En,
            Imm => ID_EX_imm,
            OUT_EN => ID_EX_OUT_En,
            CLR => '0',
            PCPlus4 => ID_EX_PCPlus4,
            WB_Waddr_Sel => ID_EX_Waddr_Sel,
            WB_Wdata_Sel => ID_EX_Wdata_Sel,

            MemRead_Out => EX_MEM_Mem_Read_En,
            MEM_OP_Out => EX_MEM_Mem_Op,
            MEM_SEL_Out => EX_MEM_Mem_Addr_Sel,
            MEM_R_Out => open,
            ALURes_Out => EX_MEM_ALU_result,
            Raddr1_Out => EX_MEM_Rsrc1,
            Raddr2_Out => EX_MEM_Rsrc2,
            Rdst_Out => EX_MEM_Rdst,
            PCPlus4_Out => EX_MEM_PCPlus4,
            PCSRC_Out => open,
            Stack_en_Out => EX_MEM_Stack_En,
            Stack_inc_Out => EX_MEM_Stack_Inc,
            Stack_dec_Out => EX_MEM_Stack_Dec,
            BR_ADDR_Out => EX_MEM_BR_ADDR,
            Rdata1_Out => EX_MEM_Rdata1,
            Rdata2_Out => EX_MEM_Rdata2,
            Mem_Wdata_Sel_Out => EX_MEM_Mem_Wdata_Sel,
            WE1_Out => EX_MEM_WE1,
            WE2_Out => EX_MEM_WE2,
            MEM_W_Out => EX_MEM_Mem_Write_En,
            IN_Port_Out => open,
            Imm_Out => EX_MEM_imm,
            OUT_EN_Out => EX_MEM_OUT_En,
            WB_Waddr_Sel_Out => EX_MEM_Waddr_Sel,
            WB_Wdata_Sel_out => EX_MEM_Wdata_Sel
        );

    EX_MEM_RegWrite <= EX_MEM_WE1;

    -- ====== MEMORY ======

    -- Stack Pointer
   -- SP_enable <= EX_MEM_Stack_En;

STACK_inst: entity work.STACK
    Port Map(
        clk => clk,
        reset => reset,
        SP_enable => EX_MEM_Stack_En,
        SP_INC => EX_MEM_Stack_Inc,
        SP_DEC => EX_MEM_Stack_Dec,
        SP_out => SP_value
    );

    -- Memory Address Mux
    process(EX_MEM_Mem_Addr_Sel, EX_MEM_ALU_result, SP_value, PC_value)
    begin
        case EX_MEM_Mem_Addr_Sel is
            when "00" =>   Mem_Addr <= PC_value;
            when "01" =>   Mem_Addr <= EX_MEM_ALU_result;
            when "10" =>   Mem_Addr <= SP_value;
            when others => Mem_Addr <= PC_value;
        end case;
    end process;

    -- Memory Write Data Mux
    process(EX_MEM_Mem_Wdata_Sel, EX_MEM_Rdata1, EX_MEM_Rdata2, EX_MEM_PCPlus4)
    begin
        case EX_MEM_Mem_Wdata_Sel is
            when "00" =>   Mem_Write_Data <= EX_MEM_Rdata1;
            when "01" =>   Mem_Write_Data <= EX_MEM_Rdata2;
            when "10" =>   Mem_Write_Data <= EX_MEM_PCPlus4;
            when others => Mem_Write_Data <= EX_MEM_Rdata1;
        end case;
    end process;

    -- ====== MEM/WB PIPELINE REGISTER ======

    M_W_Register_inst: entity work.M_W_Register
        Port Map(
            CLK => clk,
            RST => reset,
            EN => '1',
            ALURes => EX_MEM_ALU_result,
            Raddr1 => EX_MEM_Rsrc1,
            Raddr2 => EX_MEM_Rsrc2,
            Rdst => EX_MEM_Rdst,
            Rdata1 => EX_MEM_Rdata1,
            Rdata2 => EX_MEM_Rdata2,
            WE1 => EX_MEM_WE1,
            WE2 => EX_MEM_WE2,
            IN_Port => '0',
            RT_ADDR => EX_MEM_PCPlus4,
            LD_DATA => Mem_Read_Data,
            Imm => EX_MEM_imm,
            OUT_EN => EX_MEM_OUT_En,
            CLR => '0',
            WB_Waddr_Sel => EX_MEM_Waddr_Sel,
            WB_Wdata_Sel => EX_MEM_Wdata_Sel,

            ALURes_Out => MEM_WB_ALU_result,
            Raddr1_Out => MEM_WB_Rsrc1,
            Raddr2_Out => MEM_WB_Rsrc2,
            Rdst_Out => MEM_WB_Rdst,
            RT_ADDR_Out => open,
            Rdata1_Out => MEM_WB_Rdata1,
            Rdata2_Out => open,
            WE1_Out => MEM_WB_WE1,
            WE2_Out => MEM_WB_WE2,
            IN_Port_Out => open,
            LD_DATA_Out => MEM_WB_Mem_Data,
            Imm_Out => MEM_WB_imm,
            OUT_EN_Out => MEM_WB_OUT_En,
            WB_Waddr_Sel_Out => MEM_WB_Waddr_Sel,
            WB_Wdata_Sel_Out => MEM_WB_Wdata_Sel
        );

    MEM_WB_RegWrite <= MEM_WB_WE1;

    -- ====== WRITE BACK ======

    -- 000: ALURes, 001: Rdata1, 010: Rdata2, 011: IMM, 100: ALURes, 101: LD_Data, 110: IN, 111: N/A
    -- Write Back Data Mux
    process(MEM_WB_Wdata_Sel, MEM_WB_ALU_result, MEM_WB_Rdata1, MEM_WB_Mem_Data,
            MEM_WB_imm, IN_PORT, MEM_WB_IN_PORT)
    begin
        case MEM_WB_Wdata_Sel is
            when "000" =>   Reg_Wdata1 <= MEM_WB_ALU_result;
            when "001" =>   Reg_Wdata1 <= MEM_WB_Rdata1;
            when "010" =>   Reg_Wdata1 <= (others => '0');
            when "011" =>   Reg_Wdata1 <= MEM_WB_imm;
            when "100" =>   Reg_Wdata1 <= MEM_WB_ALU_result;
            when "101" =>   Reg_Wdata1 <= MEM_WB_Mem_Data;
            when "110" =>   Reg_Wdata1 <= IN_PORT;
            when others =>  Reg_Wdata1 <= MEM_WB_ALU_result;
        end case;
    end process;

    -- Write Back Address Mux
    process(MEM_WB_Waddr_Sel, MEM_WB_Rdst, MEM_WB_Rsrc1, MEM_WB_Rsrc2)
    begin
        case MEM_WB_Waddr_Sel is
            when "00" =>   Reg_Waddr1 <= MEM_WB_Rdst;
            when "01" =>   Reg_Waddr1 <= MEM_WB_Rsrc1;
            when "10" =>   Reg_Waddr1 <= MEM_WB_Rsrc2;
            when others => Reg_Waddr1 <= MEM_WB_Rdst;
        end case;
    end process;

    -- Write Enable signals
    Reg_WE1 <= MEM_WB_WE1;
    Reg_WE2 <= MEM_WB_WE2;
    Reg_Waddr2 <= (others => '0');
    Reg_Wdata2 <= (others => '0');

    -- Output Port
    process(clk, reset)
    begin
        if reset = '1' then
            OUT_PORT <= (others => '0');
        elsif rising_edge(clk) then
            if MEM_WB_OUT_En = '1' then
                OUT_PORT <= MEM_WB_Rdata1;
            end if;
        end if;
    end process;

    -- PC Write Enable
    PC_we <= '1' when PCsrc = '1' and branch_taken = '1' else '0';

    -- Flush IF/ID on branch
    --IF_ID_Flush <= '0';
    --IF_ID_Flush <= '1' when (PCsrc = '1' and branch_taken = '1') else '0';

END processor_arch;
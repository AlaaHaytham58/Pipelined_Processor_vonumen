LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY Control_Unit IS
	PORT(	
            --Inputs
            clk,rst : IN std_logic;
            opcode: IN std_logic_vector(7 downto 0);
            HW_INT: IN std_logic;
            SW_INT: IN std_logic;

            -- Rdst vs Rsrc mux selector
            Raddr_Sel: OUT STD_LOGIC; -- 0: Rsrc, 1: Rdst

            --Execute Signals
            RTI,Branch: OUT std_logic;
            Int_Jump_Sel: OUT std_logic;                -- 0 : IMM, 1: INTERRUPT
            Int_Idx : OUT STD_LOGIC_VECTOR(1 downto 0); -- 00: N/A, 01: 1, 10: 2, 11: 3
            J_Type: OUT STD_LOGIC_VECTOR(1 downto 0);   -- 00: Z, 01: N, 10: C, 11: 1
            ALU_A, ALU_B: OUT STD_LOGIC;                -- 0 : Rdata1/Rdata2, 1: Rdata2/Imm
            ALU_Op: OUT STD_LOGIC_VECTOR(2 downto 0);   -- REFER TO THE TABLE IN THE REPORT
            CCR_En: OUT STD_LOGIC;

            --Memory Signals
            Mem_Write_En, Mem_Read_En,Stack_En, PCsrc: OUT std_logic;
            Stack_Inc: OUT std_logic;                        -- 0: +4, 1: -4
            Mem_Op: OUT std_logic;
            Mem_Addr_Sel: OUT STD_LOGIC_VECTOR(1 downto 0);  -- 00: PC 01: ALURes 10: SP  
            Mem_Write_Sel: OUT STD_LOGIC_VECTOR(1 downto 0); -- 00: Rdata1 01: Rdata2 10: PCPlus4
            
            --Write Back Signals
            WE1, WE2: OUT std_logic;

            -- 00: Rdst, 01: Raddr1, 10: Raddr2, 11: ALURes
            WB_Wadrr_Sel: OUT STD_LOGIC_VECTOR(1 downto 0); 
            OUT_En : OUT STD_LOGIC;

             -- 000: ALURes, 001: Rdata1, 010: Rdata2, 011: IMM, 100: ALURes, 101: LD_Data, 110: IN, 111: N/A
            WB_Wdata_Sel: OUT STD_LOGIC_VECTOR(2 downto 0); 

            -- HLT
            HLT : OUT STD_LOGIC
        );
END Control_Unit;

ARCHITECTURE Control_Unit_arch OF Control_Unit IS
BEGIN
    process(clk, rst) begin
        -- Default Values
        Raddr_Sel <= '0';

        (RTI, Branch) <= "00";
        (Int_Idx, Int_Jump_Sel,J_Type) <= "000000";
        (ALU_A, ALU_B) <= "00";
        ALU_Op <= "00";
        CCR_En <= '0';

        (Mem_Write_En, Mem_Read_En,Stack_En, PCsrc) <= "0000";
        (Stack_Inc, Mem_Op) <= "00";
        Mem_Addr_Sel <= "00";
        Mem_Write_Sel <= "00";

        (WE1, WE2) <= "00";
        WB_Wadrr_Sel <= "00";    
        WB_Wdata_Sel <= "000";
        OUT_en <= '0';     

        HLT <= '0';
        if (CLK'event and CLK = '1' and rst = '0') then
            -- Higher priority to HW interrupt
            if (HW_INT = '1') then
                Int_Jump_Sel <= '1'; 
                Int_Idx <= "01";
            else 
                -- First 4 bits are fixed
                Mem_Op <= opcode(7);
                PCsrc  <= opcode(6);
                CCR_En <= opcode(5);
                WE1    <= opcode(4);

                -- Decode based on operation type
                case(opcode(7 downto 6)) is
                    -- ALU and Rtype operations
                    when "00" =>
                        -- ALU operations
                        if (CCR_En) then
                            -- Set opcode
                            ALU_Op <= opcode(2 downto 0);

                            -- One operand operations read from Rdst otherwise from Rsrc
                            Raddr_Sel <= '1' when opcode(2) = '1' else '0';

                            -- IADD takes immediate  in B, otherwise, rsrc2
                            ALU_B <= '1' when opcode(2 downto 0) = "101" else '0';
                        else
                        -- Rtype operations
                            HLT <= '1' when opcode(2 downto 0) = "001";
                            
                            -- Read Rsrc for move otherwise read Rdst (or don't care for operations that don't use rdata1)
                            Raddr_Sel <= '0' when opcode(2 downto 0) = "011" else '1';
                            
                            -- Write in Rdst for operations with Write back
                            WB_Wadrr_Sel <= "00";

                            -- For writing to OUT port in write operations
                            OUT_En <= '1' when opcode(2 downto 0) = "010";

                            -- To write back data for Swap
                            WE2 <= '1' when opcode(2 downto 0) = "101";
                            
                            -- WB data selection: Imm in the case of LDM, IN for IN instruction, Rdata2 for swap ,Rdata1 otherwise
                            WB_Wdata_Sel <= "011" when opcode(2 downto 0) = "110" else
                                            "111" when opcode(2 downto 0) = "001" else
                                            "010" when opcode(2 downto 0) = "101" else
                                            "001";
                        end if;    

                    -- Branch Operations                       
                    when "01" =>
                        J_Type <= opcode(1 downto 0);
                        Branch <= '1';
                    -- Memory Operations
                    when "10" =>
                        -- Choose ALURes or SP
                        Mem_Addr_Sel <= opcode(2 downto 1);

                        -- Enable MemWrite for push and std
                        Mem_Write_En <= opcode(0);

                        -- Enable MemRead for op and ldd
                        Mem_Read_En <= not opcode(0);

                        -- Enable SP for push pop
                        Stack_En <= opcode(1);

                        -- Choose increment or decrement SP
                        Stack_Inc <= opcode(0);

                        -- for load and store, ALU operands are rsrc2, Imm
                        ALU_A <= '1';
                        ALU_B <= '1';

                        -- to add offset and rsrc2 for load and store
                        ALU_OP <= "001";

                        -- to write back LD_Data for pop and ldd
                        WB_Wdata_Sel <= "101";

                    -- Branch with memory operations
                    when "11" =>
                        -- Branch during Execute in Call and INT
                        branch <= opcode(0);

                        -- Branching is always unconditional
                        J_Type <= "11";
                        
                        -- Choose intterupt or immediate for call/int (don't care otherwise)
                        Int_Jump_Sel <= opcode(1);

                        -- Choose the address that the interrupt jumps to (don't care if operation is not INT)
                        Int_Idx <= "10" when SW_INT = '0' else "11";
                        
                        -- Enable MemWrite for call, int
                        Mem_Write_En <= opcode(0);

                        -- Enable MemRead for op and ldd
                        Mem_Read_En <= not opcode(0);

                        -- Enable SP for push pop
                        Stack_En <= opcode(1);

                        -- Choose increment or decrement SP
                        Stack_Inc <= opcode(0);

                end case;
            end if;
        end if;
    end process;

END Control_Unit_arch;